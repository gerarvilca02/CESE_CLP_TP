library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package coeffs_pkg is
  constant TAPS : integer := 64;
  subtype coeff_t is signed(15 downto 0);
  type coeff_arr_t is array (0 to TAPS-1) of coeff_t;
  type coeff_bank_t is array (0 to 3) of coeff_arr_t;
  constant COEFFS : coeff_bank_t := (
    0 => (
      to_signed(37, 16), to_signed(40, 16), to_signed(46, 16), to_signed(55, 16), to_signed(68, 16), to_signed(83, 16), to_signed(102, 16), to_signed(126, 16), to_signed(153, 16), to_signed(184, 16), to_signed(219, 16), to_signed(257, 16), to_signed(300, 16), to_signed(345, 16), to_signed(393, 16), to_signed(444, 16), to_signed(496, 16), to_signed(550, 16), to_signed(604, 16), to_signed(658, 16), to_signed(712, 16), to_signed(764, 16), to_signed(814, 16), to_signed(861, 16), to_signed(905, 16), to_signed(945, 16), to_signed(981, 16), to_signed(1011, 16), to_signed(1036, 16), to_signed(1055, 16), to_signed(1067, 16), to_signed(1074, 16), to_signed(1074, 16), to_signed(1067, 16), to_signed(1055, 16), to_signed(1036, 16), to_signed(1011, 16), to_signed(981, 16), to_signed(945, 16), to_signed(905, 16), to_signed(861, 16), to_signed(814, 16), to_signed(764, 16), to_signed(712, 16), to_signed(658, 16), to_signed(604, 16), to_signed(550, 16), to_signed(496, 16), to_signed(444, 16), to_signed(393, 16), to_signed(345, 16), to_signed(300, 16), to_signed(257, 16), to_signed(219, 16), to_signed(184, 16), to_signed(153, 16), to_signed(126, 16), to_signed(102, 16), to_signed(83, 16), to_signed(68, 16), to_signed(55, 16), to_signed(46, 16), to_signed(40, 16), to_signed(37, 16)
    ),
    1 => (
      to_signed(-23, 16), to_signed(-22, 16), to_signed(-22, 16), to_signed(-22, 16), to_signed(-21, 16), to_signed(-18, 16), to_signed(-13, 16), to_signed(-6, 16), to_signed(7, 16), to_signed(24, 16), to_signed(48, 16), to_signed(78, 16), to_signed(116, 16), to_signed(163, 16), to_signed(217, 16), to_signed(280, 16), to_signed(351, 16), to_signed(429, 16), to_signed(513, 16), to_signed(602, 16), to_signed(696, 16), to_signed(791, 16), to_signed(886, 16), to_signed(979, 16), to_signed(1069, 16), to_signed(1153, 16), to_signed(1229, 16), to_signed(1295, 16), to_signed(1351, 16), to_signed(1393, 16), to_signed(1422, 16), to_signed(1437, 16), to_signed(1437, 16), to_signed(1422, 16), to_signed(1393, 16), to_signed(1351, 16), to_signed(1295, 16), to_signed(1229, 16), to_signed(1153, 16), to_signed(1069, 16), to_signed(979, 16), to_signed(886, 16), to_signed(791, 16), to_signed(696, 16), to_signed(602, 16), to_signed(513, 16), to_signed(429, 16), to_signed(351, 16), to_signed(280, 16), to_signed(217, 16), to_signed(163, 16), to_signed(116, 16), to_signed(78, 16), to_signed(48, 16), to_signed(24, 16), to_signed(7, 16), to_signed(-6, 16), to_signed(-13, 16), to_signed(-18, 16), to_signed(-21, 16), to_signed(-22, 16), to_signed(-22, 16), to_signed(-22, 16), to_signed(-23, 16)
    ),
    2 => (
      to_signed(26, 16), to_signed(25, 16), to_signed(14, 16), to_signed(-7, 16), to_signed(-33, 16), to_signed(-53, 16), to_signed(-54, 16), to_signed(-26, 16), to_signed(31, 16), to_signed(97, 16), to_signed(140, 16), to_signed(126, 16), to_signed(39, 16), to_signed(-103, 16), to_signed(-246, 16), to_signed(-313, 16), to_signed(-244, 16), to_signed(-28, 16), to_signed(275, 16), to_signed(542, 16), to_signed(626, 16), to_signed(424, 16), to_signed(-58, 16), to_signed(-682, 16), to_signed(-1195, 16), to_signed(-1303, 16), to_signed(-781, 16), to_signed(431, 16), to_signed(2176, 16), to_signed(4099, 16), to_signed(5745, 16), to_signed(6694, 16), to_signed(6694, 16), to_signed(5745, 16), to_signed(4099, 16), to_signed(2176, 16), to_signed(431, 16), to_signed(-781, 16), to_signed(-1303, 16), to_signed(-1195, 16), to_signed(-682, 16), to_signed(-58, 16), to_signed(424, 16), to_signed(626, 16), to_signed(542, 16), to_signed(275, 16), to_signed(-28, 16), to_signed(-244, 16), to_signed(-313, 16), to_signed(-246, 16), to_signed(-103, 16), to_signed(39, 16), to_signed(126, 16), to_signed(140, 16), to_signed(97, 16), to_signed(31, 16), to_signed(-26, 16), to_signed(-54, 16), to_signed(-53, 16), to_signed(-33, 16), to_signed(-7, 16), to_signed(14, 16), to_signed(25, 16), to_signed(26, 16)
    ),
    3 => (
      to_signed(-10, 16), to_signed(22, 16), to_signed(25, 16), to_signed(-14, 16), to_signed(-44, 16), to_signed(-7, 16), to_signed(60, 16), to_signed(49, 16), to_signed(-59, 16), to_signed(-108, 16), to_signed(18, 16), to_signed(166, 16), to_signed(76, 16), to_signed(-186, 16), to_signed(-217, 16), to_signed(122, 16), to_signed(368, 16), to_signed(56, 16), to_signed(-458, 16), to_signed(-348, 16), to_signed(402, 16), to_signed(706, 16), to_signed(-116, 16), to_signed(-1027, 16), to_signed(-467, 16), to_signed(1154, 16), to_signed(1402, 16), to_signed(-846, 16), to_signed(-2871, 16), to_signed(-536, 16), to_signed(6387, 16), to_signed(12683, 16), to_signed(12683, 16), to_signed(6387, 16), to_signed(-536, 16), to_signed(-2871, 16), to_signed(-846, 16), to_signed(1402, 16), to_signed(1154, 16), to_signed(-467, 16), to_signed(-1027, 16), to_signed(-116, 16), to_signed(706, 16), to_signed(402, 16), to_signed(-348, 16), to_signed(-458, 16), to_signed(56, 16), to_signed(368, 16), to_signed(122, 16), to_signed(-217, 16), to_signed(-186, 16), to_signed(76, 16), to_signed(166, 16), to_signed(18, 16), to_signed(-108, 16), to_signed(-59, 16), to_signed(49, 16), to_signed(60, 16), to_signed(-7, 16), to_signed(-44, 16), to_signed(-14, 16), to_signed(25, 16), to_signed(22, 16), to_signed(-10, 16)
    )
  );
end package coeffs_pkg;